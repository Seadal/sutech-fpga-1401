library IEEE;
use IEEE.Std_logic_1164.all;
use IEEE.Numeric_Std.all;

entity tb is

end entity;


architecture of tb is

  component WS

	Port 
		(
		temp, light, clock, reset : in std_logic;
	        moist : in std_logic_vector (2 downto 0);
		myState : out std_logic_vector(1 downto 0);
		mySeg : out std_logic_vector(6 downto 0);
		moistOut : out std_logic_vector (2 downto 0);
		tempOut : out std_logic;
		lightOut : out std_logic
		);
 end component;

	 signal temp, light, clock, reset : in std_logic;
	 signal moist : in std_logic_vector (2 downto 0);
	 signal myState : out std_logic_vector(1 downto 0);
	 signal mySeg : out std_logic_vector(6 downto 0);
	 signal moistOut : out std_logic_vector (2 downto 0);
	 signal tempOut : out std_logic;
	 signal lightOut : out std_logic

	constat cp: time := 100 ns;
	signal stop: boolean;

begin

porting : WS port map 	
	(
		temp => temp,
		light => light,
		clock => clock,
		reset => reset,
		moist => moist,
		myState => myState,
		mySeg => mySeg,
		moistOut => moistOut,
		tempOut=> tempOut,
		lightOut => lightOut
	);
ex: process

  begin

    temp <= '0';
    light <= '0';
    moist <= "110";
    wait for cp;
    temp <= '1';
    light <= '1';
    moist <= "001";
    wait for cp;
    TEMP_IN <= '0';
    LIGHT_IN <= '0';
    moist <= "101";
    wait for cp;
    temp <= '0';
    light <= '0';
    moist <= "011";
    wait for cp;
    temp <= '0';
    light <= '0';
    moist <= "111";
    wait for cp;
    temp <= '1';
    light <= '1';
    moist <= "010";
    wait for cp;
    temp <= '1';
    light <= '1';
    moist <= "011";
    wait for cp;
    temp <= '1';
    light <= '1';
    moist <= "010";
    wait for cp;


    STOP <= true;
    wait;
  end process;

  clocking: process
  begin
    while not stop loop
      clock <= '0', '1' after cp / 2;
      wait for cp;
    end loop;
    wait;
  end process;

end;


