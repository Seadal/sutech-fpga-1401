LIBRARY ieee;
USE ieee.std_logic_1164.all;

--...................................................................................--

entity seg is
	Port (
		display : in std_logic_vector ( 1 downto 0);
		ssd: out std_logic_vector (6 downto 0)
	      );
END seg;

--...................................................................................--

architecture Behavioral of seg is
	begin
		ssd <= "1001000" when display = "01" 
		else
			"1111110";
end architecture;
--...................................................................................--